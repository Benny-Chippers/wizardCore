module vga_control (

);

endmodule
