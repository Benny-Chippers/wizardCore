module id_immGen (
   i_instr,
   o_imm
);
  // I/O
  input logic [31:0] i_instr;
  output logic [31:0] o_imm;

  always_comb begin
    unique case (i_instr[6:0])
      7'b0010011: begin
        // I-Type Instruction (OP IMM)
        o_imm = {{20{i_instr[31]}}, i_instr[31:20]};
      end

      7'b0000011: begin
        // I-Type Instruction (LOAD)
        o_imm = {{20{i_instr[31]}}, i_instr[31:20]};
      end

      7'b1100111: begin
        // I-Type Instruction (JALR)
        o_imm = {{20{i_instr[31]}}, i_instr[31:20]};
      end

      7'b0100011: begin
        // S-Type Instruction (STORE)
        o_imm = {{20{i_instr[31]}}, i_instr[31:25], i_instr[11:7]};
      end

      7'b01100011: begin
        // B-Type Instruction (Branch)
        o_imm = {{19{i_instr[31]}}, i_instr[31], i_instr[7], i_instr[30:25], i_instr[11:8], 1'b0};
      end

      7'b0110111: begin
        // U-Type Instruction (Load upper immediate)
        o_imm = {i_instr[31:12], 12'b0};
      end

      7'b0010111: begin
        // U-Type Instruction (Add upper immediate to PC)
        o_imm = {i_instr[31:12], 12'b0};
      end
      7'b1101111: begin
        // J-Type Instruction (Jump and link)
        o_imm = {{11{i_instr[31]}}, i_instr[31], i_instr[19:12], i_instr[20], i_instr[30:21], 1'b0};
      end

      default: begin
        // R-Type Instruction (NOP)
        if(i_instr[0] == 1) begin
          o_imm = 32'b0;
        end else begin
          o_imm = i_instr;
        end

      end
    endcase
  end

endmodule : id_immGen
