module vga_frame (

);

endmodule
